package riscv_32i_config_pkg;
  parameter int unsigned DATA_MEM_DEPTH = 1024;
endpackage
