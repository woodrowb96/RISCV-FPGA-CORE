module alu(
  input logic [3:0] alu_op,

  input logic [31:0] in_a,
  input logic [31:0] in_b,

  output logic [31:0] result,
  output logic zero
);

endmodule
